----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:38:16 04/08/2014 
-- Design Name: 
-- Module Name:    memoriaRAM_I - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity memoriaRAM_I is port (
		  CLK : in std_logic;
		  ADDR : in std_logic_vector (31 downto 0); --Dir 
        Din : in std_logic_vector (31 downto 0);--entrada de datos para el puerto de escritura
        WE : in std_logic;		-- write enable	
		  RE : in std_logic;		-- read enable		  
		  Dout : out std_logic_vector (31 downto 0));
end memoriaRAM_I;

architecture Behavioral of memoriaRAM_I is
type RamType is array(0 to 127) of std_logic_vector(31 downto 0);

--TEST 1 ( ejemplo proporcionado en el material necesita datos1)
signal RAM : RamType := (  			X"10210003", X"1021003E", X"1021005D", X"1021006C", X"08010000", X"04212000", X"04842000", X"04844000",  -- word 0,1,2,3,4,5,6,7
									X"05088000", X"06003000", X"08040004", X"08C20000", X"10A80008", X"08C20000", X"08C20004", X"06063000", --word 8,9,...
									X"04252800", X"1000FFFB", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 16,...
									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",--word 40,...
									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
									X"08010000", X"0C017008", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",--word 72,...
									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
									X"08020104", X"0C027004", X"08020108", X"08420000", X"0C027004", X"20000000", X"00000000", X"00000000", --word 96,...
									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
									X"0802010C", X"0C027004", X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
--TEST 2 (ESCRITURA LIMPIA Y SUCIA necesita datos 1)
-- C�DIGO EN ENSAMBLADOR
--	beq R1, R1, INI;
--	beq R1, R1, RTI;
--	beq R1, R1, RT_Abort;
--	beq R1, R1, RT_UNDEF;
--	lw R1, 0(R0)					fallo ----- tag = 0 ----- set = 0 ----- via = 0
--	add R4, R1, R1
-- 	sw R4, 0(R0)					acierto ----- via = 0	
--	sw R4, 100(R0)					fallo ----- tag = 4 ----- set = 0 ----- via = 1
--	sw R0, 80(R0)					fallo ----- tag = 2 ----- set = 0 ----- via = 0
--	sw R0, 0(R0)					fallo ----- tag = 0 ----- set = 0 ----- via = 1
--	sw R6, 0(R6)					acierto ----- via = 1	
--	add R4, R4, R4
--	add R8, R4, R4
--	add R16, R8, R8
--	add R6, R16, R0
--	lw R4, 4(R0)					acierto ----- via = 1
--buc	sw R6, 0(R6)					fallo ----- tag = 0 ----- set = 1 ----- via = 0
--	sw R6, 104(R6)					fallo ----- tag = 4 ----- set = 1 ----- via = 1
--	sw R8, 84(R6)					fallo ----- tag = 2 ----- set = 1 ----- via = 0
--	sw R8, 4(R6)					fallo ----- tag = 0 ----- set = 1 ----- via = 1
--	add R6, R16, R6					por cada iteraci�n del bucle se avanza un conjunto y al avanzar mucho el 
--	add R5, R1, R5					programa acabar� cambiando los tags, estos son hasta llenar las 2 v�as de cach�. 
-- 	beq R0, R0, buc
--signal RAM : RamType := (  			X"10210003", X"1021003E", X"1021005D", X"1021006C", X"08010000", X"04212000", X"0C040000", X"0C040100",  -- word 0,1,2,3,4,5,6,7
--									X"0C000080", X"0C000000", X"00000000", X"0CC60000",X"04842000", X"04844000", X"05088000", X"06003000",--word 8,9,...
--									X"08040004", X"0CC60000", X"0CC60104", X"0CC80084", X"0CC80004", X"06063000", X"04252800", X"1000FFF9", --word 16,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",--word 40,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
--									X"08010000", X"0C017008", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",--word 72,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--									X"08020104", X"0C027004", X"08020108", X"08420000", X"0C027004", X"20000000", X"00000000", X"00000000", --word 96,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--									X"0802010C", X"0C027004", X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
--									
			

--TEST 3 (ESCRITURAS Y LECTURA EN SCRACH, necesita datos 2)
-- C�DIGO EN ENSAMBLADOR
--	beq R1, R1, INI;
--	beq R1, R1, RTI;
--	beq R1, R1, RT_Abort;
--	beq R1, R1, RT_UNDEF;
--	lw R1, 0(R0)					fallo ----- tag = 0 ----- set = 0 ----- via = 0
--	lw R2, 4(R0)					acierto ----- via = 0
--	lw R4, 8(R0)					acierto ----- via = 0
--buc	lw R3, 0(R2)					lectura de la scratch
--	add R3, R1, R3
--	add R2, R4, R2
--	sw R3, 0(R2)					escritura en la scratch
--	beq R0, R0, buc
--signal RAM : RamType := (  			X"10210003", X"1021003E", X"1021005D", X"1021006C",  X"08010000", X"08020004", X"08040008", X"08430000",   -- word 0,1,2,3,4,5,6,7
--									X"04611800", X"04441000", X"0C430000", X"1000FFFB", X"0C040080", X"08070090", X"08C20000", X"10A80008", --word 8,9,...
--									X"08C20000", X"08C20004", X"06063000", X"04252800", X"1000FFFB", X"00000000", X"00000000", X"00000000", --word 16,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",--word 40,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
--									X"08010000", X"0C017008", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",--word 72,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--									X"08020104", X"0C027004", X"08020108", X"08420000", X"0C027004", X"20000000", X"00000000", X"00000000", --word 96,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--									X"0802010C", X"0C027004", X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
--

--TEST 4 (PRUEBA 3 ERRORES)
-- C�DIGO EN ENSAMBLADOR
--	beq R1, R1, INI;
--	beq R1, R1, RTI;
--	beq R1, R1, RT_Abort;
--	beq R1, R1, RT_UNDEF;
--buc	lw R1, 111(R0)					unaligned
--	add R4, R1, R1
--	lw R1, 2110(R0)					direcci�n no detectada por la memoria
--	add R16, R8, R8
--	add R6, R16, R0
--	lw R2, 108(R0)
--	sw R3, 0(R2)					escritura en registro de lectura
--	beq R0, R0, buc
--signal RAM : RamType := (  			X"10210003", X"1021003E", X"1021005D", X"1021006C", X"08010111", X"04212000", X"04842000", X"08012110",  -- word 0,1,2,3,4,5,6,7
--									X"05088000", X"06003000", X"08020108", X"0C430000", X"1000FFF7", X"00000000", X"00000000", X"00000000", --word 8,9,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 16,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",--word 40,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
--									X"08010000", X"0C017008", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",--word 72,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--									X"08020104", X"0C027004", X"08037004", X"08020108", X"08420000", X"0C027004", X"0C087004", X"20000000", --word 96,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--									X"0802010C", X"0C027004", X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
--
--TEST 5 (COMPLETO necesita datos 2)
-- C�DIGO EN ENSAMBLADOR
--	beq R1, R1, INI;
--	beq R1, R1, RTI;
--	beq R1, R1, RT_Abort;
--	beq R1, R1, RT_UNDEF;
--	lw R1, 111(R0)						unaligned
--	lw R1, 0(R0)						fallo ----- tag = 0 ----- set = 0 ----- via = 0	
--	add R4, R1, R1						
--	add R4, R4, R4
--	lw R3, 4(R0)						acierto ----- via = 0
--	lw, R8, 4(R3)						load en la scratch
--	add R16, R8, R8
--	sw R16,4(R3)						store en la scratch
--	add R6, R16, R6
-- buc	sw R6, 0(R6)						fallo ----- tag = 0 ----- set = 1 ----- via = 0	
--	sw R6, 104(R6)						fallo ----- tag = 4 ----- set = 1 ----- via = 1
--	lw R10, 84(R6)						fallo ----- tag = 2 ----- set = 1 ----- via = 0
--	sw R8,4(R6)						fallo ----- tag = 0 ----- set = 1 ----- via = 1
--	add R6, R16, R6						por cada iteraci�n del bucle se avanza un conjunto y al avanzar mucho el 
--	add R5, R1, R5 						programa acabar� cambiando los tags, estos son hasta llenar las 2 v�as 
-- 	beq R0, R0, buc						de cach�. 

--signal RAM : RamType := (  			X"10210003", X"1021003E", X"1021005D", X"1021006C", X"08010111", X"08010000", X"04212000", X"04842000",  -- word 0,1,2,3,4,5,6,7
--									X"08030004", X"08680004", X"05088000", X"0C700004", X"06063000", X"0CC60000", X"0CC60104", X"08CA0084",--word 8,9,...
--									X"0CC80004", X"06063000",X"04252800", X"1000FFF9", X"0CC80004", X"06063000",X"04252800", X"1000FFF9", --word 16,17,...
--									X"1000FFF9", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 24,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 32,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",--word 40,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",
--									X"08010000", X"0C017008", X"20000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 64,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000",--word 72,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 80,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 88,...
--									X"08020104", X"0C027004", X"08020108", X"08420000", X"0C027004", X"20000000", X"00000000", X"00000000", --word 96,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 104,...
--									X"0802010C", X"0C027004", X"1000FFFF", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", --word 112,...
--									X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000", X"00000000");--word 120,...
--											
signal dir_7:  std_logic_vector(6 downto 0); 
begin
 
 dir_7 <= ADDR(8 downto 2); -- como la memoria es de 128 plalabras no usamos la direcci�n completa sino s�lo 7 bits. Como se direccionan los bytes, pero damos palabras no usamos los 2 bits menos significativos
 process (CLK)
    begin
        if (CLK'event and CLK = '1') then
            if (WE = '1') then -- s�lo se escribe si WE vale 1
                RAM(conv_integer(dir_7)) <= Din;
            end if;
        end if;
    end process;

    Dout <= RAM(conv_integer(dir_7)) when (RE='1') else "00000000000000000000000000000000"; --s�lo se lee si RE vale 1

end Behavioral;


